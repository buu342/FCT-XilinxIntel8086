--  C:\DOCUMENTS AND SETTINGS\SL2ALUNO\DESKTOP\NOSSO\TF2\CONTROLADOR.vhd
--  VHDL code created by Xilinx's StateCAD 9.2i
--  Fri Jun 15 00:48:33 2018

--  This VHDL code (for use with IEEE compliant tools) was generated using: 
--  binary encoded state assignment with structured code format.
--  Minimization is enabled,  implied else is enabled, 
--  and outputs are manually optimized.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SHELL_CONTROLADOR IS
	PORT (CLK,Flags0,Flags1,Flags2,Flags3,Flags4,Flags5,Flags6,Flags7,INTR,OP0,
		OP1,OP2,OP3,OP4,OP5,OP6,OP7,RESET: IN std_logic;
		DSP,EIO,ERAM,FETCH1,FETCH2,INTA,IPC,ISP,ITMP,LDTMP,nRW,RA,RB,RBus,RD,RDADD,
			RDNOT,RDXOR,RF,RIR,RMAR,RPC,RSignals,RSP,RTMP,WA,WB,WC,WD,WF,WIR,WMAR,WPC,WSP
			,WTMP,ZPC : OUT std_logic);
END;

ARCHITECTURE BEHAVIOR OF SHELL_CONTROLADOR IS
	SIGNAL sreg : std_logic_vector (6 DOWNTO 0);
	SIGNAL next_sreg : std_logic_vector (6 DOWNTO 0);
	CONSTANT CALL_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="0000000";
	CONSTANT CALL_ADDR_2 : std_logic_vector (6 DOWNTO 0) :="0000001";
	CONSTANT CALL_ADDR_3 : std_logic_vector (6 DOWNTO 0) :="0000010";
	CONSTANT CALL_ADDR_4 : std_logic_vector (6 DOWNTO 0) :="0000011";
	CONSTANT IN_C_D_1 : std_logic_vector (6 DOWNTO 0) :="0000100";
	CONSTANT IN_C_D_2 : std_logic_vector (6 DOWNTO 0) :="0000101";
	CONSTANT INT_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="0000110";
	CONSTANT INT_ADDR_2 : std_logic_vector (6 DOWNTO 0) :="0000111";
	CONSTANT INT_ADDR_3 : std_logic_vector (6 DOWNTO 0) :="0001000";
	CONSTANT INT_ADDR_4 : std_logic_vector (6 DOWNTO 0) :="0001001";
	CONSTANT INT_ADDR_5 : std_logic_vector (6 DOWNTO 0) :="0001010";
	CONSTANT INT_ADDR_6 : std_logic_vector (6 DOWNTO 0) :="0001011";
	CONSTANT INT_ADDR_7 : std_logic_vector (6 DOWNTO 0) :="0001100";
	CONSTANT INTR1 : std_logic_vector (6 DOWNTO 0) :="0001101";
	CONSTANT INTR2 : std_logic_vector (6 DOWNTO 0) :="0001110";
	CONSTANT INTR3 : std_logic_vector (6 DOWNTO 0) :="0001111";
	CONSTANT INTR4 : std_logic_vector (6 DOWNTO 0) :="0010000";
	CONSTANT INTR5 : std_logic_vector (6 DOWNTO 0) :="0010001";
	CONSTANT IRET_1 : std_logic_vector (6 DOWNTO 0) :="0010010";
	CONSTANT IRET_2 : std_logic_vector (6 DOWNTO 0) :="0010011";
	CONSTANT IRET_3 : std_logic_vector (6 DOWNTO 0) :="0010100";
	CONSTANT IRET_4 : std_logic_vector (6 DOWNTO 0) :="0010101";
	CONSTANT IRET_5 : std_logic_vector (6 DOWNTO 0) :="0010110";
	CONSTANT JMP_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="0010111";
	CONSTANT JMP_ADDR_2 : std_logic_vector (6 DOWNTO 0) :="0011000";
	CONSTANT JNZ_2_E_1 : std_logic_vector (6 DOWNTO 0) :="0011001";
	CONSTANT JNZ_2_F_1 : std_logic_vector (6 DOWNTO 0) :="0011010";
	CONSTANT JNZ_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="0011011";
	CONSTANT MOV_A_B : std_logic_vector (6 DOWNTO 0) :="0011100";
	CONSTANT MOV_A_B_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="0011101";
	CONSTANT MOV_A_B_ADDR_2 : std_logic_vector (6 DOWNTO 0) :="0011110";
	CONSTANT MOV_A_B_ADDR_3 : std_logic_vector (6 DOWNTO 0) :="0011111";
	CONSTANT MOV_A_B_ADDR_4 : std_logic_vector (6 DOWNTO 0) :="0100000";
	CONSTANT MOV_A_B_ADDR_5 : std_logic_vector (6 DOWNTO 0) :="0100001";
	CONSTANT MOV_A_B_ADDR_6 : std_logic_vector (6 DOWNTO 0) :="0100010";
	CONSTANT MOV_A_BYTE_1 : std_logic_vector (6 DOWNTO 0) :="0100011";
	CONSTANT MOV_A_BYTE_2 : std_logic_vector (6 DOWNTO 0) :="0100100";
	CONSTANT MOV_A_IBI_1 : std_logic_vector (6 DOWNTO 0) :="0100101";
	CONSTANT MOV_A_IBI_2 : std_logic_vector (6 DOWNTO 0) :="0100110";
	CONSTANT MOV_ADDR_A_1 : std_logic_vector (6 DOWNTO 0) :="0100111";
	CONSTANT MOV_ADDR_A_2 : std_logic_vector (6 DOWNTO 0) :="0101000";
	CONSTANT MOV_ADDR_A_3 : std_logic_vector (6 DOWNTO 0) :="0101001";
	CONSTANT MOV_ADDR_A_4 : std_logic_vector (6 DOWNTO 0) :="0101010";
	CONSTANT MOV_B_BYTE_1 : std_logic_vector (6 DOWNTO 0) :="0101011";
	CONSTANT MOV_B_BYTE_2 : std_logic_vector (6 DOWNTO 0) :="0101100";
	CONSTANT MOV_D_A : std_logic_vector (6 DOWNTO 0) :="0101101";
	CONSTANT MOVE_SP_BYTE_1 : std_logic_vector (6 DOWNTO 0) :="0101110";
	CONSTANT MOVE_SP_BYTE_2 : std_logic_vector (6 DOWNTO 0) :="0101111";
	CONSTANT OUT_D_B_1 : std_logic_vector (6 DOWNTO 0) :="0110000";
	CONSTANT OUT_D_B_2 : std_logic_vector (6 DOWNTO 0) :="0110001";
	CONSTANT POP_B_1 : std_logic_vector (6 DOWNTO 0) :="0110010";
	CONSTANT POP_B_2 : std_logic_vector (6 DOWNTO 0) :="0110011";
	CONSTANT POP_B_3 : std_logic_vector (6 DOWNTO 0) :="0110100";
	CONSTANT PUSH_A_1 : std_logic_vector (6 DOWNTO 0) :="0110101";
	CONSTANT PUSH_A_2 : std_logic_vector (6 DOWNTO 0) :="0110110";
	CONSTANT PUSHFLAGS_1 : std_logic_vector (6 DOWNTO 0) :="0110111";
	CONSTANT PUSHFLAGS_2 : std_logic_vector (6 DOWNTO 0) :="0111000";
	CONSTANT RET_1 : std_logic_vector (6 DOWNTO 0) :="0111001";
	CONSTANT RET_2 : std_logic_vector (6 DOWNTO 0) :="0111010";
	CONSTANT RET_3 : std_logic_vector (6 DOWNTO 0) :="0111011";
	CONSTANT STATE0 : std_logic_vector (6 DOWNTO 0) :="0111100";
	CONSTANT STATE1 : std_logic_vector (6 DOWNTO 0) :="0111101";
	CONSTANT STATE2 : std_logic_vector (6 DOWNTO 0) :="0111110";
	CONSTANT STOP : std_logic_vector (6 DOWNTO 0) :="0111111";
	CONSTANT SUB_A_ADDR_1 : std_logic_vector (6 DOWNTO 0) :="1000000";
	CONSTANT SUB_A_ADDR_2 : std_logic_vector (6 DOWNTO 0) :="1000001";
	CONSTANT SUB_A_ADDR_3 : std_logic_vector (6 DOWNTO 0) :="1000010";
	CONSTANT SUB_A_ADDR_4 : std_logic_vector (6 DOWNTO 0) :="1000011";
	CONSTANT SUB_A_ADDR_5 : std_logic_vector (6 DOWNTO 0) :="1000100";
	CONSTANT SUB_A_ADDR_6 : std_logic_vector (6 DOWNTO 0) :="1000101";
	CONSTANT SUB_A_ADDR_7 : std_logic_vector (6 DOWNTO 0) :="1000110";
	CONSTANT XOR_B_A_1 : std_logic_vector (6 DOWNTO 0) :="1000111";
	CONSTANT XOR_B_A_2 : std_logic_vector (6 DOWNTO 0) :="1001000";
	CONSTANT XOR_B_A_3 : std_logic_vector (6 DOWNTO 0) :="1001001";

BEGIN
	PROCESS (CLK, RESET, next_sreg)
	BEGIN
		IF ( RESET='1' ) THEN
			sreg <= STATE0;
		ELSIF CLK='0' AND CLK'event THEN
			sreg <= next_sreg;
		END IF;
	END PROCESS;

	PROCESS (sreg,Flags4,INTR,OP0,OP1,OP2,OP3,OP4,OP5,OP6,OP7)
	BEGIN
		DSP <= '0'; EIO <= '0'; ERAM <= '0'; FETCH1 <= '0'; FETCH2 <= '0'; INTA <= 
			'0'; IPC <= '0'; ISP <= '0'; ITMP <= '0'; LDTMP <= '0'; nRW <= '0'; RA <= 
			'0'; RB <= '0'; RBus <= '0'; RD <= '0'; RDADD <= '0'; RDNOT <= '0'; RDXOR <= 
			'0'; RF <= '0'; RIR <= '0'; RMAR <= '0'; RPC <= '0'; RSignals <= '0'; RSP <= 
			'0'; RTMP <= '0'; WA <= '0'; WB <= '0'; WC <= '0'; WD <= '0'; WF <= '0'; WIR 
			<= '0'; WMAR <= '0'; WPC <= '0'; WSP <= '0'; WTMP <= '0'; ZPC <= '0'; 

		next_sreg<=CALL_ADDR_1;

		CASE sreg IS
			WHEN CALL_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				LDTMP<='1';
				WTMP<='1';
				next_sreg<=CALL_ADDR_2;
			WHEN CALL_ADDR_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WPC<='1';
				ITMP<='1';
				next_sreg<=CALL_ADDR_3;
			WHEN CALL_ADDR_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=CALL_ADDR_4;
			WHEN CALL_ADDR_4 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				nRW<='1';
				DSP<='1';
				RTMP<='1';
				next_sreg<=STATE1;
			WHEN IN_C_D_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RD<='1';
				WMAR<='1';
				next_sreg<=IN_C_D_2;
			WHEN IN_C_D_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				DSP<='0';
				RMAR<='1';
				WC<='1';
				EIO<='1';
				next_sreg<=STATE1;
			WHEN INT_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=INT_ADDR_2;
			WHEN INT_ADDR_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				IPC<='1';
				WIR<='1';
				next_sreg<=INT_ADDR_3;
			WHEN INT_ADDR_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=INT_ADDR_4;
			WHEN INT_ADDR_4 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				RF<='1';
				nRW<='1';
				DSP<='1';
				next_sreg<=INT_ADDR_5;
			WHEN INT_ADDR_5 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=INT_ADDR_6;
			WHEN INT_ADDR_6 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				nRW<='1';
				RPC<='1';
				next_sreg<=INT_ADDR_7;
			WHEN INT_ADDR_7 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='1';
				RIR<='1';
				WPC<='1';
				next_sreg<=STATE1;
			WHEN INTR1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=INTR2;
			WHEN INTR2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				nRW<='1';
				RF<='1';
				DSP<='1';
				next_sreg<=INTR3;
			WHEN INTR3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=INTR4;
			WHEN INTR4 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				nRW<='1';
				RPC<='1';
				DSP<='1';
				next_sreg<=INTR5;
			WHEN INTR5 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				WPC<='1';
				INTA<='1';
				next_sreg<=STATE1;
			WHEN IRET_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				ISP<='1';
				next_sreg<=IRET_2;
			WHEN IRET_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=IRET_3;
			WHEN IRET_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WPC<='1';
				ISP<='1';
				next_sreg<=IRET_4;
			WHEN IRET_4 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=IRET_5;
			WHEN IRET_5 =>
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WF<='1';
				RBus<='1';
				next_sreg<=STATE1;
			WHEN JMP_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=JMP_ADDR_2;
			WHEN JMP_ADDR_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WPC<='1';
				next_sreg<=STATE1;
			WHEN JNZ_2_E_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				IPC<='1';
				next_sreg<=STATE1;
			WHEN JNZ_2_F_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WPC<='1';
				next_sreg<=STATE1;
			WHEN JNZ_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				IF ( Flags4='0' ) THEN
					next_sreg<=JNZ_2_F_1;
				 ELSE
					next_sreg<=JNZ_2_E_1;
				END IF;
			WHEN MOV_A_B =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RB<='1';
				WA<='1';
				next_sreg<=STATE1;
			WHEN MOV_A_B_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=MOV_A_B_ADDR_2;
			WHEN MOV_A_B_ADDR_2 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				LDTMP<='1';
				WTMP<='1';
				IPC<='1';
				next_sreg<=MOV_A_B_ADDR_3;
			WHEN MOV_A_B_ADDR_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RTMP<='1';
				WMAR<='1';
				next_sreg<=MOV_A_B_ADDR_4;
			WHEN MOV_A_B_ADDR_4 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				LDTMP<='1';
				WTMP<='1';
				next_sreg<=MOV_A_B_ADDR_5;
			WHEN MOV_A_B_ADDR_5 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RD<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RB<='1';
				RDADD<='1';
				WTMP<='1';
				RSignals<='1';
				WF<='1';
				next_sreg<=MOV_A_B_ADDR_6;
			WHEN MOV_A_B_ADDR_6 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RTMP<='1';
				WA<='1';
				next_sreg<=STATE1;
			WHEN MOV_A_BYTE_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=MOV_A_BYTE_2;
			WHEN MOV_A_BYTE_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WA<='1';
				IPC<='1';
				next_sreg<=STATE1;
			WHEN MOV_A_IBI_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RB<='1';
				WMAR<='1';
				next_sreg<=MOV_A_IBI_2;
			WHEN MOV_A_IBI_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				ERAM<='1';
				WA<='1';
				RMAR<='1';
				next_sreg<=STATE1;
			WHEN MOV_ADDR_A_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=MOV_ADDR_A_2;
			WHEN MOV_ADDR_A_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WIR<='1';
				IPC<='1';
				next_sreg<=MOV_ADDR_A_3;
			WHEN MOV_ADDR_A_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RIR<='1';
				WMAR<='1';
				next_sreg<=MOV_ADDR_A_4;
			WHEN MOV_ADDR_A_4 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				RA<='1';
				nRW<='1';
				next_sreg<=STATE1;
			WHEN MOV_B_BYTE_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=MOV_B_BYTE_2;
			WHEN MOV_B_BYTE_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WB<='1';
				IPC<='1';
				next_sreg<=STATE1;
			WHEN MOV_D_A =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RA<='1';
				WD<='1';
				next_sreg<=STATE1;
			WHEN MOVE_SP_BYTE_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=MOVE_SP_BYTE_2;
			WHEN MOVE_SP_BYTE_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				IPC<='1';
				WSP<='1';
				next_sreg<=STATE1;
			WHEN OUT_D_B_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RD<='1';
				WMAR<='1';
				next_sreg<=OUT_D_B_2;
			WHEN OUT_D_B_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				DSP<='0';
				RMAR<='1';
				RB<='1';
				EIO<='1';
				nRW<='1';
				next_sreg<=STATE1;
			WHEN POP_B_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				ISP<='1';
				next_sreg<=POP_B_2;
			WHEN POP_B_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=POP_B_3;
			WHEN POP_B_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WB<='1';
				next_sreg<=STATE1;
			WHEN PUSH_A_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=PUSH_A_2;
			WHEN PUSH_A_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				nRW<='1';
				RA<='1';
				DSP<='1';
				next_sreg<=STATE1;
			WHEN PUSHFLAGS_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=PUSHFLAGS_2;
			WHEN PUSHFLAGS_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				RMAR<='1';
				ERAM<='1';
				RF<='1';
				nRW<='1';
				DSP<='1';
				next_sreg<=STATE1;
			WHEN RET_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				ISP<='1';
				next_sreg<=RET_2;
			WHEN RET_2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RSP<='1';
				WMAR<='1';
				next_sreg<=RET_3;
			WHEN RET_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WPC<='1';
				next_sreg<=STATE1;
			WHEN STATE0 =>
				RBus<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				ZPC<='1';
				next_sreg<=STATE1;
			WHEN STATE1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				FETCH1<='1';
				IF ( INTR='1' ) THEN
					next_sreg<=INTR1;
				 ELSE
					next_sreg<=STATE2;
				END IF;
			WHEN STATE2 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WIR<='1';
				IPC<='1';
				FETCH2<='1';
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='1' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=MOV_A_B;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='0' 
					AND OP1='1' AND OP0='1' ) THEN
					next_sreg<=MOV_D_A;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='0' 
					AND OP1='1' AND OP0='0' ) THEN
					next_sreg<=JNZ_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='0' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=IRET_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='0' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=INT_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='1' 
					AND OP1='1' AND OP0='0' ) THEN
					next_sreg<=CALL_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='1' 
					AND OP1='1' AND OP0='0' ) THEN
					next_sreg<=MOV_A_IBI_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='0' 
					AND OP1='1' AND OP0='0' ) THEN
					next_sreg<=MOV_A_B_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='1' 
					AND OP1='1' AND OP0='1' ) THEN
					next_sreg<=STOP;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='0' 
					AND OP1='1' AND OP0='1' ) THEN
					next_sreg<=XOR_B_A_1;
				END IF;
				IF ( OP7='1' ) OR ( OP6='1' ) OR ( OP5='1' ) OR ( OP3='1' AND OP4='1' ) 
					OR ( OP1='1' AND OP2='1' AND OP4='1' ) THEN
					next_sreg<=STATE1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='0' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=MOV_A_BYTE_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='0' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=SUB_A_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='1' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=MOV_B_BYTE_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='0' AND OP2='1' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=MOV_ADDR_A_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='0' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=IN_C_D_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='0' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=OUT_D_B_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='0' 
					AND OP1='1' AND OP0='0' ) THEN
					next_sreg<=PUSH_A_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='0' 
					AND OP1='1' AND OP0='1' ) THEN
					next_sreg<=POP_B_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='1' 
					AND OP1='0' AND OP0='0' ) THEN
					next_sreg<=JMP_ADDR_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='1' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=RET_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='0' AND OP3='1' AND OP2='1' 
					AND OP1='1' AND OP0='1' ) THEN
					next_sreg<=MOVE_SP_BYTE_1;
				END IF;
				IF ( OP7='0' AND OP6='0' AND OP5='0' AND OP4='1' AND OP3='0' AND OP2='1' 
					AND OP1='0' AND OP0='1' ) THEN
					next_sreg<=PUSHFLAGS_1;
				END IF;
			WHEN STOP =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				next_sreg<=STOP;
			WHEN SUB_A_ADDR_1 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RPC<='1';
				WMAR<='1';
				next_sreg<=SUB_A_ADDR_2;
			WHEN SUB_A_ADDR_2 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WTMP<='1';
				LDTMP<='1';
				next_sreg<=SUB_A_ADDR_3;
			WHEN SUB_A_ADDR_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RTMP<='1';
				WMAR<='1';
				next_sreg<=SUB_A_ADDR_4;
			WHEN SUB_A_ADDR_4 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				EIO<='0';
				DSP<='0';
				RMAR<='1';
				ERAM<='1';
				WTMP<='1';
				RDNOT<='1';
				next_sreg<=SUB_A_ADDR_5;
			WHEN SUB_A_ADDR_5 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				ITMP<='1';
				next_sreg<=SUB_A_ADDR_6;
			WHEN SUB_A_ADDR_6 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RD<='0';
				RB<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RA<='1';
				RDADD<='1';
				WTMP<='1';
				RSignals<='1';
				WF<='1';
				next_sreg<=SUB_A_ADDR_7;
			WHEN SUB_A_ADDR_7 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RTMP<='1';
				WA<='1';
				IPC<='1';
				next_sreg<=STATE1;
			WHEN XOR_B_A_1 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RA<='0';
				nRW<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RB<='1';
				WTMP<='1';
				LDTMP<='1';
				next_sreg<=XOR_B_A_2;
			WHEN XOR_B_A_2 =>
				RBus<='0';
				ZPC<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WD<='0';
				WC<='0';
				WB<='0';
				WA<='0';
				RTMP<='0';
				RSP<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RA<='1';
				RDXOR<='1';
				WTMP<='1';
				RSignals<='1';
				WF<='1';
				next_sreg<=XOR_B_A_3;
			WHEN XOR_B_A_3 =>
				RBus<='0';
				ZPC<='0';
				WTMP<='0';
				WSP<='0';
				WPC<='0';
				WMAR<='0';
				WIR<='0';
				WF<='0';
				WD<='0';
				WC<='0';
				WA<='0';
				RSP<='0';
				RSignals<='0';
				RPC<='0';
				RMAR<='0';
				RIR<='0';
				RF<='0';
				RDXOR<='0';
				RDNOT<='0';
				RDADD<='0';
				RD<='0';
				RB<='0';
				RA<='0';
				nRW<='0';
				LDTMP<='0';
				ITMP<='0';
				ISP<='0';
				IPC<='0';
				INTA<='0';
				FETCH2<='0';
				FETCH1<='0';
				ERAM<='0';
				EIO<='0';
				DSP<='0';
				RTMP<='1';
				WB<='1';
				next_sreg<=STATE1;
			WHEN OTHERS =>
		END CASE;
	END PROCESS;
END BEHAVIOR;

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CONTROLADOR IS
	PORT (FLAGS : IN std_logic_vector (7 DOWNTO 0);
		OP : IN std_logic_vector (7 DOWNTO 0);
		CLK,INTR,RESET: IN std_logic;
		DSP,EIO,ERAM,FETCH1,FETCH2,INTA,IPC,ISP,ITMP,LDTMP,nRW,RA,RB,RBus,RD,RDADD,
			RDNOT,RDXOR,RF,RIR,RMAR,RPC,RSignals,RSP,RTMP,WA,WB,WC,WD,WF,WIR,WMAR,WPC,WSP
			,WTMP,ZPC : OUT std_logic);
END;

ARCHITECTURE BEHAVIOR OF CONTROLADOR IS
	COMPONENT SHELL_CONTROLADOR
		PORT (CLK,Flags0,Flags1,Flags2,Flags3,Flags4,Flags5,Flags6,Flags7,INTR,OP0,
			OP1,OP2,OP3,OP4,OP5,OP6,OP7,RESET: IN std_logic;
			DSP,EIO,ERAM,FETCH1,FETCH2,INTA,IPC,ISP,ITMP,LDTMP,nRW,RA,RB,RBus,RD,RDADD
				,RDNOT,RDXOR,RF,RIR,RMAR,RPC,RSignals,RSP,RTMP,WA,WB,WC,WD,WF,WIR,WMAR,WPC,
				WSP,WTMP,ZPC : OUT std_logic);
	END COMPONENT;
BEGIN
	SHELL1_CONTROLADOR : SHELL_CONTROLADOR PORT MAP (CLK=>CLK,Flags0=>FLAGS(0),
		Flags1=>FLAGS(1),Flags2=>FLAGS(2),Flags3=>FLAGS(3),Flags4=>FLAGS(4),Flags5=>
		FLAGS(5),Flags6=>FLAGS(6),Flags7=>FLAGS(7),INTR=>INTR,OP0=>OP(0),OP1=>OP(1),
		OP2=>OP(2),OP3=>OP(3),OP4=>OP(4),OP5=>OP(5),OP6=>OP(6),OP7=>OP(7),RESET=>
		RESET,DSP=>DSP,EIO=>EIO,ERAM=>ERAM,FETCH1=>FETCH1,FETCH2=>FETCH2,INTA=>INTA,
		IPC=>IPC,ISP=>ISP,ITMP=>ITMP,LDTMP=>LDTMP,nRW=>nRW,RA=>RA,RB=>RB,RBus=>RBus,
		RD=>RD,RDADD=>RDADD,RDNOT=>RDNOT,RDXOR=>RDXOR,RF=>RF,RIR=>RIR,RMAR=>RMAR,RPC
		=>RPC,RSignals=>RSignals,RSP=>RSP,RTMP=>RTMP,WA=>WA,WB=>WB,WC=>WC,WD=>WD,WF=>
		WF,WIR=>WIR,WMAR=>WMAR,WPC=>WPC,WSP=>WSP,WTMP=>WTMP,ZPC=>ZPC);
END BEHAVIOR;
